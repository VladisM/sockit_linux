library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SoCkit_Linux is port(
	OSC_50_B8A									  : in 	 std_logic;												-- clock
	
	memory_mem_a                    		  : out   std_logic_vector(14 downto 0);              -- mem_a
	memory_mem_ba                   		  : out   std_logic_vector(2 downto 0);               -- mem_ba
	memory_mem_ck                   		  : out   std_logic;                                  -- mem_ck
	memory_mem_ck_n                 		  : out   std_logic;                                  -- mem_ck_n
	memory_mem_cke                  		  : out   std_logic;                                  -- mem_cke
	memory_mem_cs_n                		  : out   std_logic;                                  -- mem_cs_n
	memory_mem_ras_n                		  : out   std_logic;                                  -- mem_ras_n
	memory_mem_cas_n                		  : out   std_logic;                                  -- mem_cas_n
	memory_mem_we_n                 		  : out   std_logic;                                  -- mem_we_n
	memory_mem_reset_n              		  : out   std_logic;                                  -- mem_reset_n
	memory_mem_dq                   		  : inout std_logic_vector(31 downto 0);					-- mem_dq
	memory_mem_dqs                 		  : inout std_logic_vector(3 downto 0);               -- mem_dqs
	memory_mem_dqs_n               		  : inout std_logic_vector(3 downto 0);               -- mem_dqs_n
	memory_mem_odt                  		  : out   std_logic;                                  -- mem_odt
	memory_mem_dm                   		  : out   std_logic_vector(3 downto 0);               -- mem_dm
	memory_oct_rzqin                		  : in    std_logic;                                  -- oct_rzqin
	
	hps_0_hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                  -- hps_io_emac1_inst_TX_CLK
	hps_0_hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                  -- hps_io_emac1_inst_TXD0
	hps_0_hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                  -- hps_io_emac1_inst_TXD1
	hps_0_hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                  -- hps_io_emac1_inst_TXD2
	hps_0_hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                  -- hps_io_emac1_inst_TXD3
	hps_0_hps_io_hps_io_emac1_inst_RXD0   : in    std_logic;             							-- hps_io_emac1_inst_RXD0
	hps_0_hps_io_hps_io_emac1_inst_MDIO   : inout std_logic;           								-- hps_io_emac1_inst_MDIO
	hps_0_hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                  -- hps_io_emac1_inst_MDC
	hps_0_hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic;             							-- hps_io_emac1_inst_RX_CTL
	hps_0_hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                  -- hps_io_emac1_inst_TX_CTL
	hps_0_hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic;             							-- hps_io_emac1_inst_RX_CLK
	hps_0_hps_io_hps_io_emac1_inst_RXD1   : in    std_logic;             							-- hps_io_emac1_inst_RXD1
	hps_0_hps_io_hps_io_emac1_inst_RXD2   : in    std_logic;             							-- hps_io_emac1_inst_RXD2
	hps_0_hps_io_hps_io_emac1_inst_RXD3   : in    std_logic;             							-- hps_io_emac1_inst_RXD3

	hps_0_hps_io_hps_io_sdio_inst_CMD     : inout std_logic;         									-- hps_io_sdio_inst_CMD
	hps_0_hps_io_hps_io_sdio_inst_D0      : inout std_logic;           							   -- hps_io_sdio_inst_D0
	hps_0_hps_io_hps_io_sdio_inst_D1      : inout std_logic;            								-- hps_io_sdio_inst_D1
	hps_0_hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                  -- hps_io_sdio_inst_CLK
	hps_0_hps_io_hps_io_sdio_inst_D2      : inout std_logic;                             		-- hps_io_sdio_inst_D2
	hps_0_hps_io_hps_io_sdio_inst_D3      : inout std_logic;   											-- hps_io_sdio_inst_D3
			
	hps_0_hps_io_hps_io_uart0_inst_RX     : in    std_logic;                     					-- hps_io_uart0_inst_RX
	hps_0_hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                  -- hps_io_uart0_inst_TX

	LED											  : out std_logic_vector(3 downto 0);						-- leds 
	KEY											  : in std_logic_vector(3 downto 0);						-- push buttons
	SW												  : in std_logic_vector(3 downto 0));						-- switchs 
end entity SoCkit_Linux;
		
architecture main of SoCkit_Linux is		
	component SoC is port (
		memory_mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
		memory_mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
		memory_mem_ck                   : out   std_logic;                                        -- mem_ck
		memory_mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
		memory_mem_cke                  : out   std_logic;                                        -- mem_cke
		memory_mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
		memory_mem_ras_n                : out   std_logic;                                        -- mem_ras_n
		memory_mem_cas_n                : out   std_logic;                                        -- mem_cas_n
		memory_mem_we_n                 : out   std_logic;                                        -- mem_we_n
		memory_mem_reset_n              : out   std_logic;                                        -- mem_reset_n
		memory_mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
		memory_mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
		memory_mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
		memory_mem_odt                  : out   std_logic;                                        -- mem_odt
		memory_mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
		memory_oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin

		hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3

		hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3

		hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX

		reset_reset_n                   : in    std_logic                     := 'X';             -- reset_n
		clk_clk                         : in    std_logic                     := 'X';             -- clk

		sw_export                       : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
		led_export                      : out   std_logic_vector(7 downto 0));                    -- export
	end component SoC;

	signal led_signal: std_logic_vector(7 downto 0);
	signal sw_signal: std_logic_vector(7 downto 0);
	
begin

	sw_signal(3 downto 0) <= KEY;
	sw_signal(7 downto 4) <= SW;
	LED <= led_signal(3 downto 0);

	u0 : component SoC
		port map (
			memory_mem_a                    => memory_mem_a,                          --                  memory.mem_a
			memory_mem_ba                   => memory_mem_ba,                         --                        .mem_ba
			memory_mem_ck                   => memory_mem_ck,                         --                        .mem_ck
			memory_mem_ck_n                 => memory_mem_ck_n,                       --                        .mem_ck_n
			memory_mem_cke                  => memory_mem_cke,                        --                        .mem_cke
			memory_mem_cs_n                 => memory_mem_cs_n,                       --                        .mem_cs_n
			memory_mem_ras_n                => memory_mem_ras_n,                		  --                        .mem_ras_n
			memory_mem_cas_n                => memory_mem_cas_n,            		     --                        .mem_cas_n
			memory_mem_we_n                 => memory_mem_we_n,              		     --                        .mem_we_n
			memory_mem_reset_n              => memory_mem_reset_n,           			  --                        .mem_reset_n
			memory_mem_dq                   => memory_mem_dq,                 		  --                        .mem_dq
			memory_mem_dqs                  => memory_mem_dqs,                		  --                        .mem_dqs
			memory_mem_dqs_n                => memory_mem_dqs_n,               		  --                        .mem_dqs_n
			memory_mem_odt                  => memory_mem_odt,                  		  --                        .mem_odt
			memory_mem_dm                   => memory_mem_dm,                   		  --                        .mem_dm
			memory_oct_rzqin                => memory_oct_rzqin,                		  --                        .oct_rzqin
			
			hps_io_hps_io_emac1_inst_TX_CLK => hps_0_hps_io_hps_io_emac1_inst_TX_CLK, --                  hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_hps_io_emac1_inst_TXD0   => hps_0_hps_io_hps_io_emac1_inst_TXD0,   --                        .hps_io_emac1_inst_TXD0
			hps_io_hps_io_emac1_inst_TXD1   => hps_0_hps_io_hps_io_emac1_inst_TXD1,   --                        .hps_io_emac1_inst_TXD1
			hps_io_hps_io_emac1_inst_TXD2   => hps_0_hps_io_hps_io_emac1_inst_TXD2,   --                        .hps_io_emac1_inst_TXD2
			hps_io_hps_io_emac1_inst_TXD3   => hps_0_hps_io_hps_io_emac1_inst_TXD3,   --                        .hps_io_emac1_inst_TXD3
			hps_io_hps_io_emac1_inst_RXD0   => hps_0_hps_io_hps_io_emac1_inst_RXD0,   --                        .hps_io_emac1_inst_RXD0
			hps_io_hps_io_emac1_inst_MDIO   => hps_0_hps_io_hps_io_emac1_inst_MDIO,   --                        .hps_io_emac1_inst_MDIO
			hps_io_hps_io_emac1_inst_MDC    => hps_0_hps_io_hps_io_emac1_inst_MDC,    --                        .hps_io_emac1_inst_MDC
			hps_io_hps_io_emac1_inst_RX_CTL => hps_0_hps_io_hps_io_emac1_inst_RX_CTL, --                        .hps_io_emac1_inst_RX_CTL
			hps_io_hps_io_emac1_inst_TX_CTL => hps_0_hps_io_hps_io_emac1_inst_TX_CTL, --                        .hps_io_emac1_inst_TX_CTL
			hps_io_hps_io_emac1_inst_RX_CLK => hps_0_hps_io_hps_io_emac1_inst_RX_CLK, --                        .hps_io_emac1_inst_RX_CLK
			hps_io_hps_io_emac1_inst_RXD1   => hps_0_hps_io_hps_io_emac1_inst_RXD1,   --                        .hps_io_emac1_inst_RXD1
			hps_io_hps_io_emac1_inst_RXD2   => hps_0_hps_io_hps_io_emac1_inst_RXD2,   --                        .hps_io_emac1_inst_RXD2
			hps_io_hps_io_emac1_inst_RXD3   => hps_0_hps_io_hps_io_emac1_inst_RXD3,   --                        .hps_io_emac1_inst_RXD3
			
			hps_io_hps_io_sdio_inst_CMD     => hps_0_hps_io_hps_io_sdio_inst_CMD,     --                        .hps_io_sdio_inst_CMD
			hps_io_hps_io_sdio_inst_D0      => hps_0_hps_io_hps_io_sdio_inst_D0,      --                        .hps_io_sdio_inst_D0
			hps_io_hps_io_sdio_inst_D1      => hps_0_hps_io_hps_io_sdio_inst_D1,      --                        .hps_io_sdio_inst_D1
			hps_io_hps_io_sdio_inst_CLK     => hps_0_hps_io_hps_io_sdio_inst_CLK,     --                        .hps_io_sdio_inst_CLK
			hps_io_hps_io_sdio_inst_D2      => hps_0_hps_io_hps_io_sdio_inst_D2,      --                        .hps_io_sdio_inst_D2
			hps_io_hps_io_sdio_inst_D3      => hps_0_hps_io_hps_io_sdio_inst_D3,      --                        .hps_io_sdio_inst_D3
			
			hps_io_hps_io_uart0_inst_RX     => hps_0_hps_io_hps_io_uart0_inst_RX,     --                        .hps_io_uart0_inst_RX
			hps_io_hps_io_uart0_inst_TX     => hps_0_hps_io_hps_io_uart0_inst_TX,     --                        .hps_io_uart0_inst_TX

			reset_reset_n                   => '1',              						     --  					  reset.reset_n
			clk_clk                         => OSC_50_B8A,                       	  --    						 clk.clk

			sw_export                       => sw_signal,       			              --     					  sw.export
			led_export                      => led_signal 		                       --    						 led.export
		);
end architecture main;