-- soc_system.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.05.02.16:00:40

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		clk_clk                         : in    std_logic                     := '0';             --                     clk.clk
		reset_reset_n                   : in    std_logic                     := '0';             --                   reset.reset_n
		memory_mem_a                    : out   std_logic_vector(14 downto 0);                    --                  memory.mem_a
		memory_mem_ba                   : out   std_logic_vector(2 downto 0);                     --                        .mem_ba
		memory_mem_ck                   : out   std_logic;                                        --                        .mem_ck
		memory_mem_ck_n                 : out   std_logic;                                        --                        .mem_ck_n
		memory_mem_cke                  : out   std_logic;                                        --                        .mem_cke
		memory_mem_cs_n                 : out   std_logic;                                        --                        .mem_cs_n
		memory_mem_ras_n                : out   std_logic;                                        --                        .mem_ras_n
		memory_mem_cas_n                : out   std_logic;                                        --                        .mem_cas_n
		memory_mem_we_n                 : out   std_logic;                                        --                        .mem_we_n
		memory_mem_reset_n              : out   std_logic;                                        --                        .mem_reset_n
		memory_mem_dq                   : inout std_logic_vector(31 downto 0) := (others => '0'); --                        .mem_dq
		memory_mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs
		memory_mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => '0'); --                        .mem_dqs_n
		memory_mem_odt                  : out   std_logic;                                        --                        .mem_odt
		memory_mem_dm                   : out   std_logic_vector(3 downto 0);                     --                        .mem_dm
		memory_oct_rzqin                : in    std_logic                     := '0';             --                        .oct_rzqin
		hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --                  hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --                        .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --                        .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --                        .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --                        .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --                        .hps_io_emac1_inst_RXD3
		hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --                        .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --                        .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := '0';             --                        .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := '0';             --                        .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP     : out   std_logic;                                        --                        .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := '0';             --                        .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := '0';             --                        .hps_io_usb1_inst_NXT
		hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --                        .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --                        .hps_io_uart0_inst_TX
		led_external_connection_export  : out   std_logic_vector(7 downto 0);                     -- led_external_connection.export
		pb_external_connection_export   : in    std_logic_vector(7 downto 0)  := (others => '0')  --  pb_external_connection.export
	);
end entity soc_system;

architecture rtl of soc_system is
	component soc_system_hps is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                        -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component soc_system_hps;

	component soc_system_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component soc_system_led;

	component soc_system_pb is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component soc_system_pb;

	component number_generator is
		port (
			reset_in : in  std_logic                     := 'X'; -- reset_n
			clk_in   : in  std_logic                     := 'X'; -- clk
			CS       : in  std_logic                     := 'X'; -- chipselect
			OE       : in  std_logic                     := 'X'; -- read
			readdata : out std_logic_vector(31 downto 0)         -- readdata
		);
	end component number_generator;

	component altera_merlin_axi_master_ni is
		generic (
			ID_WIDTH                  : integer := 2;
			ADDR_WIDTH                : integer := 32;
			RDATA_WIDTH               : integer := 32;
			WDATA_WIDTH               : integer := 32;
			ADDR_USER_WIDTH           : integer := 5;
			DATA_USER_WIDTH           : integer := 8;
			AXI_BURST_LENGTH_WIDTH    : integer := 4;
			AXI_LOCK_WIDTH            : integer := 2;
			AXI_VERSION               : string  := "AXI3";
			WRITE_ISSUING_CAPABILITY  : integer := 16;
			READ_ISSUING_CAPABILITY   : integer := 16;
			PKT_BEGIN_BURST           : integer := 104;
			PKT_CACHE_H               : integer := 103;
			PKT_CACHE_L               : integer := 100;
			PKT_ADDR_SIDEBAND_H       : integer := 99;
			PKT_ADDR_SIDEBAND_L       : integer := 92;
			PKT_PROTECTION_H          : integer := 89;
			PKT_PROTECTION_L          : integer := 87;
			PKT_BURST_SIZE_H          : integer := 84;
			PKT_BURST_SIZE_L          : integer := 82;
			PKT_BURST_TYPE_H          : integer := 86;
			PKT_BURST_TYPE_L          : integer := 85;
			PKT_RESPONSE_STATUS_L     : integer := 106;
			PKT_RESPONSE_STATUS_H     : integer := 107;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_EXCLUSIVE       : integer := 81;
			PKT_TRANS_LOCK            : integer := 105;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 109;
			PKT_THREAD_ID_L           : integer := 108;
			PKT_QOS_L                 : integer := 110;
			PKT_QOS_H                 : integer := 113;
			PKT_DATA_SIDEBAND_H       : integer := 121;
			PKT_DATA_SIDEBAND_L       : integer := 114;
			ST_DATA_W                 : integer := 122;
			ST_CHANNEL_W              : integer := 1;
			ID                        : integer := 1
		);
		port (
			aclk                   : in  std_logic                      := 'X';             -- clk
			aresetn                : in  std_logic                      := 'X';             -- reset_n
			write_cp_valid         : out std_logic;                                         -- valid
			write_cp_data          : out std_logic_vector(110 downto 0);                    -- data
			write_cp_startofpacket : out std_logic;                                         -- startofpacket
			write_cp_endofpacket   : out std_logic;                                         -- endofpacket
			write_cp_ready         : in  std_logic                      := 'X';             -- ready
			write_rp_valid         : in  std_logic                      := 'X';             -- valid
			write_rp_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			write_rp_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			write_rp_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			write_rp_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			write_rp_ready         : out std_logic;                                         -- ready
			read_cp_valid          : out std_logic;                                         -- valid
			read_cp_data           : out std_logic_vector(110 downto 0);                    -- data
			read_cp_startofpacket  : out std_logic;                                         -- startofpacket
			read_cp_endofpacket    : out std_logic;                                         -- endofpacket
			read_cp_ready          : in  std_logic                      := 'X';             -- ready
			read_rp_valid          : in  std_logic                      := 'X';             -- valid
			read_rp_data           : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			read_rp_channel        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			read_rp_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			read_rp_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			read_rp_ready          : out std_logic;                                         -- ready
			awid                   : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			awaddr                 : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- awaddr
			awlen                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			awsize                 : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			awburst                : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			awlock                 : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			awcache                : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			awprot                 : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			awvalid                : in  std_logic                      := 'X';             -- awvalid
			awready                : out std_logic;                                         -- awready
			wid                    : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			wdata                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- wdata
			wstrb                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- wstrb
			wlast                  : in  std_logic                      := 'X';             -- wlast
			wvalid                 : in  std_logic                      := 'X';             -- wvalid
			wready                 : out std_logic;                                         -- wready
			bid                    : out std_logic_vector(11 downto 0);                     -- bid
			bresp                  : out std_logic_vector(1 downto 0);                      -- bresp
			bvalid                 : out std_logic;                                         -- bvalid
			bready                 : in  std_logic                      := 'X';             -- bready
			arid                   : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			araddr                 : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- araddr
			arlen                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			arsize                 : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			arburst                : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			arlock                 : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			arcache                : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			arprot                 : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			arvalid                : in  std_logic                      := 'X';             -- arvalid
			arready                : out std_logic;                                         -- arready
			rid                    : out std_logic_vector(11 downto 0);                     -- rid
			rdata                  : out std_logic_vector(31 downto 0);                     -- rdata
			rresp                  : out std_logic_vector(1 downto 0);                      -- rresp
			rlast                  : out std_logic;                                         -- rlast
			rvalid                 : out std_logic;                                         -- rvalid
			rready                 : in  std_logic                      := 'X';             -- rready
			awuser                 : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- awuser
			aruser                 : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- aruser
			awqos                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awqos
			arqos                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arqos
			awregion               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awregion
			arregion               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arregion
			wuser                  : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- wuser
			ruser                  : out std_logic_vector(0 downto 0);                      -- ruser
			buser                  : out std_logic_vector(0 downto 0)                       -- buser
		);
	end component altera_merlin_axi_master_ni;

	component altera_merlin_slave_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(20 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(110 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(111 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(111 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_agent;

	component soc_system_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(110 downto 0);                    -- data
			src_channel        : out std_logic_vector(2 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component soc_system_addr_router;

	component soc_system_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(110 downto 0);                    -- data
			src_channel        : out std_logic_vector(2 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component soc_system_id_router;

	component altera_merlin_traffic_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(110 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(2 downto 0);                      -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(110 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(2 downto 0);                      -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(2 downto 0)                       -- data
		);
	end component altera_merlin_traffic_limiter;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                      := 'X';             -- clk
			reset                 : in  std_logic                      := 'X';             -- reset
			sink0_valid           : in  std_logic                      := 'X';             -- valid
			sink0_data            : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                         -- ready
			source0_valid         : out std_logic;                                         -- valid
			source0_data          : out std_logic_vector(110 downto 0);                    -- data
			source0_channel       : out std_logic_vector(2 downto 0);                      -- channel
			source0_startofpacket : out std_logic;                                         -- startofpacket
			source0_endofpacket   : out std_logic;                                         -- endofpacket
			source0_ready         : in  std_logic                      := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component soc_system_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(110 downto 0);                    -- data
			src0_channel       : out std_logic_vector(2 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(110 downto 0);                    -- data
			src1_channel       : out std_logic_vector(2 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(110 downto 0);                    -- data
			src2_channel       : out std_logic_vector(2 downto 0);                      -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component soc_system_cmd_xbar_demux;

	component soc_system_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(110 downto 0);                    -- data
			src_channel         : out std_logic_vector(2 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component soc_system_cmd_xbar_mux;

	component soc_system_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(110 downto 0);                    -- data
			src0_channel       : out std_logic_vector(2 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(110 downto 0);                    -- data
			src1_channel       : out std_logic_vector(2 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component soc_system_rsp_xbar_demux;

	component soc_system_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(110 downto 0);                    -- data
			src_channel         : out std_logic_vector(2 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component soc_system_rsp_xbar_mux;

	component soc_system_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_led_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component soc_system_led_s1_translator;

	component soc_system_pb_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component soc_system_pb_s1_translator;

	component soc_system_lfsr_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component soc_system_lfsr_0_avalon_slave_0_translator;

	component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(111 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(111 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(33 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	signal led_s1_translator_avalon_anti_slave_0_writedata                                            : std_logic_vector(31 downto 0);  -- led_s1_translator:av_writedata -> led:writedata
	signal led_s1_translator_avalon_anti_slave_0_address                                              : std_logic_vector(1 downto 0);   -- led_s1_translator:av_address -> led:address
	signal led_s1_translator_avalon_anti_slave_0_chipselect                                           : std_logic;                      -- led_s1_translator:av_chipselect -> led:chipselect
	signal led_s1_translator_avalon_anti_slave_0_write                                                : std_logic;                      -- led_s1_translator:av_write -> led_s1_translator_avalon_anti_slave_0_write:in
	signal led_s1_translator_avalon_anti_slave_0_readdata                                             : std_logic_vector(31 downto 0);  -- led:readdata -> led_s1_translator:av_readdata
	signal pb_s1_translator_avalon_anti_slave_0_address                                               : std_logic_vector(1 downto 0);   -- pb_s1_translator:av_address -> pb:address
	signal pb_s1_translator_avalon_anti_slave_0_readdata                                              : std_logic_vector(31 downto 0);  -- pb:readdata -> pb_s1_translator:av_readdata
	signal lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect                            : std_logic;                      -- lfsr_0_avalon_slave_0_translator:av_chipselect -> lfsr_0:CS
	signal lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- lfsr_0_avalon_slave_0_translator:av_read -> lfsr_0:OE
	signal lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- lfsr_0:readdata -> lfsr_0_avalon_slave_0_translator:av_readdata
	signal hps_h2f_lw_axi_master_awvalid                                                              : std_logic;                      -- hps:h2f_lw_AWVALID -> hps_h2f_lw_axi_master_agent:awvalid
	signal hps_h2f_lw_axi_master_arsize                                                               : std_logic_vector(2 downto 0);   -- hps:h2f_lw_ARSIZE -> hps_h2f_lw_axi_master_agent:arsize
	signal hps_h2f_lw_axi_master_arlock                                                               : std_logic_vector(1 downto 0);   -- hps:h2f_lw_ARLOCK -> hps_h2f_lw_axi_master_agent:arlock
	signal hps_h2f_lw_axi_master_awcache                                                              : std_logic_vector(3 downto 0);   -- hps:h2f_lw_AWCACHE -> hps_h2f_lw_axi_master_agent:awcache
	signal hps_h2f_lw_axi_master_arready                                                              : std_logic;                      -- hps_h2f_lw_axi_master_agent:arready -> hps:h2f_lw_ARREADY
	signal hps_h2f_lw_axi_master_arid                                                                 : std_logic_vector(11 downto 0);  -- hps:h2f_lw_ARID -> hps_h2f_lw_axi_master_agent:arid
	signal hps_h2f_lw_axi_master_rready                                                               : std_logic;                      -- hps:h2f_lw_RREADY -> hps_h2f_lw_axi_master_agent:rready
	signal hps_h2f_lw_axi_master_bready                                                               : std_logic;                      -- hps:h2f_lw_BREADY -> hps_h2f_lw_axi_master_agent:bready
	signal hps_h2f_lw_axi_master_awsize                                                               : std_logic_vector(2 downto 0);   -- hps:h2f_lw_AWSIZE -> hps_h2f_lw_axi_master_agent:awsize
	signal hps_h2f_lw_axi_master_awprot                                                               : std_logic_vector(2 downto 0);   -- hps:h2f_lw_AWPROT -> hps_h2f_lw_axi_master_agent:awprot
	signal hps_h2f_lw_axi_master_arvalid                                                              : std_logic;                      -- hps:h2f_lw_ARVALID -> hps_h2f_lw_axi_master_agent:arvalid
	signal hps_h2f_lw_axi_master_arprot                                                               : std_logic_vector(2 downto 0);   -- hps:h2f_lw_ARPROT -> hps_h2f_lw_axi_master_agent:arprot
	signal hps_h2f_lw_axi_master_bid                                                                  : std_logic_vector(11 downto 0);  -- hps_h2f_lw_axi_master_agent:bid -> hps:h2f_lw_BID
	signal hps_h2f_lw_axi_master_arlen                                                                : std_logic_vector(3 downto 0);   -- hps:h2f_lw_ARLEN -> hps_h2f_lw_axi_master_agent:arlen
	signal hps_h2f_lw_axi_master_awready                                                              : std_logic;                      -- hps_h2f_lw_axi_master_agent:awready -> hps:h2f_lw_AWREADY
	signal hps_h2f_lw_axi_master_awid                                                                 : std_logic_vector(11 downto 0);  -- hps:h2f_lw_AWID -> hps_h2f_lw_axi_master_agent:awid
	signal hps_h2f_lw_axi_master_bvalid                                                               : std_logic;                      -- hps_h2f_lw_axi_master_agent:bvalid -> hps:h2f_lw_BVALID
	signal hps_h2f_lw_axi_master_wid                                                                  : std_logic_vector(11 downto 0);  -- hps:h2f_lw_WID -> hps_h2f_lw_axi_master_agent:wid
	signal hps_h2f_lw_axi_master_awlock                                                               : std_logic_vector(1 downto 0);   -- hps:h2f_lw_AWLOCK -> hps_h2f_lw_axi_master_agent:awlock
	signal hps_h2f_lw_axi_master_awburst                                                              : std_logic_vector(1 downto 0);   -- hps:h2f_lw_AWBURST -> hps_h2f_lw_axi_master_agent:awburst
	signal hps_h2f_lw_axi_master_bresp                                                                : std_logic_vector(1 downto 0);   -- hps_h2f_lw_axi_master_agent:bresp -> hps:h2f_lw_BRESP
	signal hps_h2f_lw_axi_master_wstrb                                                                : std_logic_vector(3 downto 0);   -- hps:h2f_lw_WSTRB -> hps_h2f_lw_axi_master_agent:wstrb
	signal hps_h2f_lw_axi_master_rvalid                                                               : std_logic;                      -- hps_h2f_lw_axi_master_agent:rvalid -> hps:h2f_lw_RVALID
	signal hps_h2f_lw_axi_master_wdata                                                                : std_logic_vector(31 downto 0);  -- hps:h2f_lw_WDATA -> hps_h2f_lw_axi_master_agent:wdata
	signal hps_h2f_lw_axi_master_wready                                                               : std_logic;                      -- hps_h2f_lw_axi_master_agent:wready -> hps:h2f_lw_WREADY
	signal hps_h2f_lw_axi_master_arburst                                                              : std_logic_vector(1 downto 0);   -- hps:h2f_lw_ARBURST -> hps_h2f_lw_axi_master_agent:arburst
	signal hps_h2f_lw_axi_master_rdata                                                                : std_logic_vector(31 downto 0);  -- hps_h2f_lw_axi_master_agent:rdata -> hps:h2f_lw_RDATA
	signal hps_h2f_lw_axi_master_araddr                                                               : std_logic_vector(20 downto 0);  -- hps:h2f_lw_ARADDR -> hps_h2f_lw_axi_master_agent:araddr
	signal hps_h2f_lw_axi_master_arcache                                                              : std_logic_vector(3 downto 0);   -- hps:h2f_lw_ARCACHE -> hps_h2f_lw_axi_master_agent:arcache
	signal hps_h2f_lw_axi_master_awlen                                                                : std_logic_vector(3 downto 0);   -- hps:h2f_lw_AWLEN -> hps_h2f_lw_axi_master_agent:awlen
	signal hps_h2f_lw_axi_master_awaddr                                                               : std_logic_vector(20 downto 0);  -- hps:h2f_lw_AWADDR -> hps_h2f_lw_axi_master_agent:awaddr
	signal hps_h2f_lw_axi_master_rid                                                                  : std_logic_vector(11 downto 0);  -- hps_h2f_lw_axi_master_agent:rid -> hps:h2f_lw_RID
	signal hps_h2f_lw_axi_master_wvalid                                                               : std_logic;                      -- hps:h2f_lw_WVALID -> hps_h2f_lw_axi_master_agent:wvalid
	signal hps_h2f_lw_axi_master_rresp                                                                : std_logic_vector(1 downto 0);   -- hps_h2f_lw_axi_master_agent:rresp -> hps:h2f_lw_RRESP
	signal hps_h2f_lw_axi_master_wlast                                                                : std_logic;                      -- hps:h2f_lw_WLAST -> hps_h2f_lw_axi_master_agent:wlast
	signal hps_h2f_lw_axi_master_rlast                                                                : std_logic;                      -- hps_h2f_lw_axi_master_agent:rlast -> hps:h2f_lw_RLAST
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                            : std_logic;                      -- led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                             : std_logic_vector(2 downto 0);   -- led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_writedata                              : std_logic_vector(31 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_address                                : std_logic_vector(20 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_write                                  : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_lock                                   : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_read                                   : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_readdata                               : std_logic_vector(31 downto 0);  -- led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                          : std_logic;                      -- led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                            : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	signal led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                             : std_logic_vector(3 downto 0);   -- led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                     : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                           : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                   : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_data                            : std_logic_vector(111 downto 0); -- led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                           : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                  : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                        : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                         : std_logic_vector(111 downto 0); -- led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                        : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                      : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                       : std_logic_vector(33 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                      : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                      : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                       : std_logic_vector(33 downto 0);  -- led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                      : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                             : std_logic;                      -- pb_s1_translator:uav_waitrequest -> pb_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                              : std_logic_vector(2 downto 0);   -- pb_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pb_s1_translator:uav_burstcount
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_writedata                               : std_logic_vector(31 downto 0);  -- pb_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pb_s1_translator:uav_writedata
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_address                                 : std_logic_vector(20 downto 0);  -- pb_s1_translator_avalon_universal_slave_0_agent:m0_address -> pb_s1_translator:uav_address
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_write                                   : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:m0_write -> pb_s1_translator:uav_write
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_lock                                    : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pb_s1_translator:uav_lock
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_read                                    : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:m0_read -> pb_s1_translator:uav_read
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                : std_logic_vector(31 downto 0);  -- pb_s1_translator:uav_readdata -> pb_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                           : std_logic;                      -- pb_s1_translator:uav_readdatavalid -> pb_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                             : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pb_s1_translator:uav_debugaccess
	signal pb_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                              : std_logic_vector(3 downto 0);   -- pb_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pb_s1_translator:uav_byteenable
	signal pb_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                      : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pb_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                            : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pb_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                    : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pb_s1_translator_avalon_universal_slave_0_agent_rf_source_data                             : std_logic_vector(111 downto 0); -- pb_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pb_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                            : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pb_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                   : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pb_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                         : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pb_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                 : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pb_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                          : std_logic_vector(111 downto 0); -- pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pb_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                         : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                       : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                        : std_logic_vector(33 downto 0);  -- pb_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                       : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pb_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                       : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pb_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                        : std_logic_vector(33 downto 0);  -- pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pb_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                       : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- lfsr_0_avalon_slave_0_translator:uav_waitrequest -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> lfsr_0_avalon_slave_0_translator:uav_burstcount
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> lfsr_0_avalon_slave_0_translator:uav_writedata
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(20 downto 0);  -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> lfsr_0_avalon_slave_0_translator:uav_address
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> lfsr_0_avalon_slave_0_translator:uav_write
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> lfsr_0_avalon_slave_0_translator:uav_lock
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> lfsr_0_avalon_slave_0_translator:uav_read
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- lfsr_0_avalon_slave_0_translator:uav_readdata -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- lfsr_0_avalon_slave_0_translator:uav_readdatavalid -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lfsr_0_avalon_slave_0_translator:uav_debugaccess
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> lfsr_0_avalon_slave_0_translator:uav_byteenable
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(111 downto 0); -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(111 downto 0); -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid       : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data        : std_logic_vector(33 downto 0);  -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready       : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal hps_h2f_lw_axi_master_agent_write_cp_endofpacket                                           : std_logic;                      -- hps_h2f_lw_axi_master_agent:write_cp_endofpacket -> addr_router:sink_endofpacket
	signal hps_h2f_lw_axi_master_agent_write_cp_valid                                                 : std_logic;                      -- hps_h2f_lw_axi_master_agent:write_cp_valid -> addr_router:sink_valid
	signal hps_h2f_lw_axi_master_agent_write_cp_startofpacket                                         : std_logic;                      -- hps_h2f_lw_axi_master_agent:write_cp_startofpacket -> addr_router:sink_startofpacket
	signal hps_h2f_lw_axi_master_agent_write_cp_data                                                  : std_logic_vector(110 downto 0); -- hps_h2f_lw_axi_master_agent:write_cp_data -> addr_router:sink_data
	signal hps_h2f_lw_axi_master_agent_write_cp_ready                                                 : std_logic;                      -- addr_router:sink_ready -> hps_h2f_lw_axi_master_agent:write_cp_ready
	signal hps_h2f_lw_axi_master_agent_read_cp_endofpacket                                            : std_logic;                      -- hps_h2f_lw_axi_master_agent:read_cp_endofpacket -> addr_router_001:sink_endofpacket
	signal hps_h2f_lw_axi_master_agent_read_cp_valid                                                  : std_logic;                      -- hps_h2f_lw_axi_master_agent:read_cp_valid -> addr_router_001:sink_valid
	signal hps_h2f_lw_axi_master_agent_read_cp_startofpacket                                          : std_logic;                      -- hps_h2f_lw_axi_master_agent:read_cp_startofpacket -> addr_router_001:sink_startofpacket
	signal hps_h2f_lw_axi_master_agent_read_cp_data                                                   : std_logic_vector(110 downto 0); -- hps_h2f_lw_axi_master_agent:read_cp_data -> addr_router_001:sink_data
	signal hps_h2f_lw_axi_master_agent_read_cp_ready                                                  : std_logic;                      -- addr_router_001:sink_ready -> hps_h2f_lw_axi_master_agent:read_cp_ready
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                            : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_valid                                  : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                          : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_data                                   : std_logic_vector(110 downto 0); -- led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal led_s1_translator_avalon_universal_slave_0_agent_rp_ready                                  : std_logic;                      -- id_router:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pb_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                             : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal pb_s1_translator_avalon_universal_slave_0_agent_rp_valid                                   : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal pb_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                           : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal pb_s1_translator_avalon_universal_slave_0_agent_rp_data                                    : std_logic_vector(110 downto 0); -- pb_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal pb_s1_translator_avalon_universal_slave_0_agent_rp_ready                                   : std_logic;                      -- id_router_001:sink_ready -> pb_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(110 downto 0); -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_002:sink_ready -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                : std_logic;                      -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                      : std_logic;                      -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                              : std_logic;                      -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                       : std_logic_vector(110 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                    : std_logic_vector(2 downto 0);   -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                      : std_logic;                      -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                : std_logic;                      -- limiter:rsp_src_endofpacket -> hps_h2f_lw_axi_master_agent:write_rp_endofpacket
	signal limiter_rsp_src_valid                                                                      : std_logic;                      -- limiter:rsp_src_valid -> hps_h2f_lw_axi_master_agent:write_rp_valid
	signal limiter_rsp_src_startofpacket                                                              : std_logic;                      -- limiter:rsp_src_startofpacket -> hps_h2f_lw_axi_master_agent:write_rp_startofpacket
	signal limiter_rsp_src_data                                                                       : std_logic_vector(110 downto 0); -- limiter:rsp_src_data -> hps_h2f_lw_axi_master_agent:write_rp_data
	signal limiter_rsp_src_channel                                                                    : std_logic_vector(2 downto 0);   -- limiter:rsp_src_channel -> hps_h2f_lw_axi_master_agent:write_rp_channel
	signal limiter_rsp_src_ready                                                                      : std_logic;                      -- hps_h2f_lw_axi_master_agent:write_rp_ready -> limiter:rsp_src_ready
	signal addr_router_001_src_endofpacket                                                            : std_logic;                      -- addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	signal addr_router_001_src_valid                                                                  : std_logic;                      -- addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	signal addr_router_001_src_startofpacket                                                          : std_logic;                      -- addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	signal addr_router_001_src_data                                                                   : std_logic_vector(110 downto 0); -- addr_router_001:src_data -> limiter_001:cmd_sink_data
	signal addr_router_001_src_channel                                                                : std_logic_vector(2 downto 0);   -- addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	signal addr_router_001_src_ready                                                                  : std_logic;                      -- limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	signal limiter_001_rsp_src_endofpacket                                                            : std_logic;                      -- limiter_001:rsp_src_endofpacket -> hps_h2f_lw_axi_master_agent:read_rp_endofpacket
	signal limiter_001_rsp_src_valid                                                                  : std_logic;                      -- limiter_001:rsp_src_valid -> hps_h2f_lw_axi_master_agent:read_rp_valid
	signal limiter_001_rsp_src_startofpacket                                                          : std_logic;                      -- limiter_001:rsp_src_startofpacket -> hps_h2f_lw_axi_master_agent:read_rp_startofpacket
	signal limiter_001_rsp_src_data                                                                   : std_logic_vector(110 downto 0); -- limiter_001:rsp_src_data -> hps_h2f_lw_axi_master_agent:read_rp_data
	signal limiter_001_rsp_src_channel                                                                : std_logic_vector(2 downto 0);   -- limiter_001:rsp_src_channel -> hps_h2f_lw_axi_master_agent:read_rp_channel
	signal limiter_001_rsp_src_ready                                                                  : std_logic;                      -- hps_h2f_lw_axi_master_agent:read_rp_ready -> limiter_001:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                          : std_logic;                      -- burst_adapter:source0_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                : std_logic;                      -- burst_adapter:source0_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                        : std_logic;                      -- burst_adapter:source0_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                 : std_logic_vector(110 downto 0); -- burst_adapter:source0_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                : std_logic;                      -- led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                              : std_logic_vector(2 downto 0);   -- burst_adapter:source0_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                      : std_logic;                      -- burst_adapter_001:source0_endofpacket -> pb_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                            : std_logic;                      -- burst_adapter_001:source0_valid -> pb_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                    : std_logic;                      -- burst_adapter_001:source0_startofpacket -> pb_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                             : std_logic_vector(110 downto 0); -- burst_adapter_001:source0_data -> pb_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                            : std_logic;                      -- pb_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                          : std_logic_vector(2 downto 0);   -- burst_adapter_001:source0_channel -> pb_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_002_source0_endofpacket                                                      : std_logic;                      -- burst_adapter_002:source0_endofpacket -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_002_source0_valid                                                            : std_logic;                      -- burst_adapter_002:source0_valid -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_002_source0_startofpacket                                                    : std_logic;                      -- burst_adapter_002:source0_startofpacket -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_002_source0_data                                                             : std_logic_vector(110 downto 0); -- burst_adapter_002:source0_data -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_002_source0_ready                                                            : std_logic;                      -- lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	signal burst_adapter_002_source0_channel                                                          : std_logic_vector(2 downto 0);   -- burst_adapter_002:source0_channel -> lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                             : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, id_router:reset, id_router_001:reset, id_router_002:reset, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lfsr_0_avalon_slave_0_translator:reset, lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, pb_s1_translator:reset, pb_s1_translator_avalon_universal_slave_0_agent:reset, pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in]
	signal hps_h2f_reset_reset                                                                        : std_logic;                      -- hps:h2f_rst_n -> hps_h2f_reset_reset:in
	signal cmd_xbar_demux_src0_endofpacket                                                            : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                  : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                          : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                   : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                : std_logic_vector(2 downto 0);   -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                  : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                            : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                  : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                          : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                   : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                : std_logic_vector(2 downto 0);   -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                  : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                            : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                  : std_logic;                      -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                          : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                   : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                : std_logic_vector(2 downto 0);   -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                  : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                              : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                      : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                               : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                            : std_logic_vector(2 downto 0);   -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                              : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                              : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                      : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                               : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                            : std_logic_vector(2 downto 0);   -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                              : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                              : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                      : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                               : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                            : std_logic_vector(2 downto 0);   -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                              : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal rsp_xbar_demux_src0_endofpacket                                                            : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                  : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                          : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                   : std_logic_vector(110 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                : std_logic_vector(2 downto 0);   -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                  : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                            : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                  : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                          : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                   : std_logic_vector(110 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                : std_logic_vector(2 downto 0);   -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                  : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                        : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                              : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                      : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                               : std_logic_vector(110 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                            : std_logic_vector(2 downto 0);   -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                              : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                        : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                              : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                      : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                               : std_logic_vector(110 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                            : std_logic_vector(2 downto 0);   -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                              : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                        : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                              : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                      : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                               : std_logic_vector(110 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                            : std_logic_vector(2 downto 0);   -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                              : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                        : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                              : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                      : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                               : std_logic_vector(110 downto 0); -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                            : std_logic_vector(2 downto 0);   -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                              : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal limiter_cmd_src_endofpacket                                                                : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                              : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                       : std_logic_vector(110 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                    : std_logic_vector(2 downto 0);   -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                      : std_logic;                      -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                               : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                     : std_logic;                      -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                             : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                      : std_logic_vector(110 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                   : std_logic_vector(2 downto 0);   -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                     : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal limiter_001_cmd_src_endofpacket                                                            : std_logic;                      -- limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal limiter_001_cmd_src_startofpacket                                                          : std_logic;                      -- limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal limiter_001_cmd_src_data                                                                   : std_logic_vector(110 downto 0); -- limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	signal limiter_001_cmd_src_channel                                                                : std_logic_vector(2 downto 0);   -- limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	signal limiter_001_cmd_src_ready                                                                  : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                           : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                 : std_logic;                      -- rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                         : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                  : std_logic_vector(110 downto 0); -- rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	signal rsp_xbar_mux_001_src_channel                                                               : std_logic_vector(2 downto 0);   -- rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	signal rsp_xbar_mux_001_src_ready                                                                 : std_logic;                      -- limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                               : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> burst_adapter:sink0_endofpacket
	signal cmd_xbar_mux_src_valid                                                                     : std_logic;                      -- cmd_xbar_mux:src_valid -> burst_adapter:sink0_valid
	signal cmd_xbar_mux_src_startofpacket                                                             : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> burst_adapter:sink0_startofpacket
	signal cmd_xbar_mux_src_data                                                                      : std_logic_vector(110 downto 0); -- cmd_xbar_mux:src_data -> burst_adapter:sink0_data
	signal cmd_xbar_mux_src_channel                                                                   : std_logic_vector(2 downto 0);   -- cmd_xbar_mux:src_channel -> burst_adapter:sink0_channel
	signal cmd_xbar_mux_src_ready                                                                     : std_logic;                      -- burst_adapter:sink0_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                  : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                        : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                         : std_logic_vector(110 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                      : std_logic_vector(2 downto 0);   -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                        : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                           : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                 : std_logic;                      -- cmd_xbar_mux_001:src_valid -> burst_adapter_001:sink0_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                         : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                  : std_logic_vector(110 downto 0); -- cmd_xbar_mux_001:src_data -> burst_adapter_001:sink0_data
	signal cmd_xbar_mux_001_src_channel                                                               : std_logic_vector(2 downto 0);   -- cmd_xbar_mux_001:src_channel -> burst_adapter_001:sink0_channel
	signal cmd_xbar_mux_001_src_ready                                                                 : std_logic;                      -- burst_adapter_001:sink0_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                              : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                    : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                            : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                     : std_logic_vector(110 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                  : std_logic_vector(2 downto 0);   -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                    : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                           : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                 : std_logic;                      -- cmd_xbar_mux_002:src_valid -> burst_adapter_002:sink0_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                         : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                  : std_logic_vector(110 downto 0); -- cmd_xbar_mux_002:src_data -> burst_adapter_002:sink0_data
	signal cmd_xbar_mux_002_src_channel                                                               : std_logic_vector(2 downto 0);   -- cmd_xbar_mux_002:src_channel -> burst_adapter_002:sink0_channel
	signal cmd_xbar_mux_002_src_ready                                                                 : std_logic;                      -- burst_adapter_002:sink0_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                              : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                    : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                            : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                     : std_logic_vector(110 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                  : std_logic_vector(2 downto 0);   -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                    : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal limiter_cmd_valid_data                                                                     : std_logic_vector(2 downto 0);   -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal limiter_001_cmd_valid_data                                                                 : std_logic_vector(2 downto 0);   -- limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	signal hps_f2h_irq0_irq                                                                           : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> hps:f2h_irq_p0
	signal hps_f2h_irq1_irq                                                                           : std_logic_vector(31 downto 0);  -- irq_mapper_001:sender_irq -> hps:f2h_irq_p1
	signal led_s1_translator_avalon_anti_slave_0_write_ports_inv                                      : std_logic;                      -- led_s1_translator_avalon_anti_slave_0_write:inv -> led:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                   : std_logic;                      -- rst_controller_reset_out_reset:inv -> [hps_h2f_lw_axi_master_agent:aresetn, led:reset_n, lfsr_0:reset_in, pb:reset_n]
	signal hps_h2f_reset_reset_ports_inv                                                              : std_logic;                      -- hps_h2f_reset_reset:inv -> rst_controller:reset_in0

begin

	hps : component soc_system_hps
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => memory_mem_a,                    --            memory.mem_a
			mem_ba                   => memory_mem_ba,                   --                  .mem_ba
			mem_ck                   => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                   --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                  --                  .mem_odt
			mem_dm                   => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK, --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,   --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,   --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,   --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,   --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,   --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,   --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,    --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL, --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL, --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK, --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,   --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,   --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,   --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,     --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,      --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,      --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,     --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,      --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,      --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,      --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,      --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,      --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,      --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,      --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,      --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,      --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,      --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,     --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,     --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,     --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,     --                  .hps_io_usb1_inst_NXT
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,     --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,     --                  .hps_io_uart0_inst_TX
			h2f_rst_n                => hps_h2f_reset_reset,             --         h2f_reset.reset_n
			h2f_lw_axi_clk           => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_h2f_lw_axi_master_awid,      -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_h2f_lw_axi_master_awaddr,    --                  .awaddr
			h2f_lw_AWLEN             => hps_h2f_lw_axi_master_awlen,     --                  .awlen
			h2f_lw_AWSIZE            => hps_h2f_lw_axi_master_awsize,    --                  .awsize
			h2f_lw_AWBURST           => hps_h2f_lw_axi_master_awburst,   --                  .awburst
			h2f_lw_AWLOCK            => hps_h2f_lw_axi_master_awlock,    --                  .awlock
			h2f_lw_AWCACHE           => hps_h2f_lw_axi_master_awcache,   --                  .awcache
			h2f_lw_AWPROT            => hps_h2f_lw_axi_master_awprot,    --                  .awprot
			h2f_lw_AWVALID           => hps_h2f_lw_axi_master_awvalid,   --                  .awvalid
			h2f_lw_AWREADY           => hps_h2f_lw_axi_master_awready,   --                  .awready
			h2f_lw_WID               => hps_h2f_lw_axi_master_wid,       --                  .wid
			h2f_lw_WDATA             => hps_h2f_lw_axi_master_wdata,     --                  .wdata
			h2f_lw_WSTRB             => hps_h2f_lw_axi_master_wstrb,     --                  .wstrb
			h2f_lw_WLAST             => hps_h2f_lw_axi_master_wlast,     --                  .wlast
			h2f_lw_WVALID            => hps_h2f_lw_axi_master_wvalid,    --                  .wvalid
			h2f_lw_WREADY            => hps_h2f_lw_axi_master_wready,    --                  .wready
			h2f_lw_BID               => hps_h2f_lw_axi_master_bid,       --                  .bid
			h2f_lw_BRESP             => hps_h2f_lw_axi_master_bresp,     --                  .bresp
			h2f_lw_BVALID            => hps_h2f_lw_axi_master_bvalid,    --                  .bvalid
			h2f_lw_BREADY            => hps_h2f_lw_axi_master_bready,    --                  .bready
			h2f_lw_ARID              => hps_h2f_lw_axi_master_arid,      --                  .arid
			h2f_lw_ARADDR            => hps_h2f_lw_axi_master_araddr,    --                  .araddr
			h2f_lw_ARLEN             => hps_h2f_lw_axi_master_arlen,     --                  .arlen
			h2f_lw_ARSIZE            => hps_h2f_lw_axi_master_arsize,    --                  .arsize
			h2f_lw_ARBURST           => hps_h2f_lw_axi_master_arburst,   --                  .arburst
			h2f_lw_ARLOCK            => hps_h2f_lw_axi_master_arlock,    --                  .arlock
			h2f_lw_ARCACHE           => hps_h2f_lw_axi_master_arcache,   --                  .arcache
			h2f_lw_ARPROT            => hps_h2f_lw_axi_master_arprot,    --                  .arprot
			h2f_lw_ARVALID           => hps_h2f_lw_axi_master_arvalid,   --                  .arvalid
			h2f_lw_ARREADY           => hps_h2f_lw_axi_master_arready,   --                  .arready
			h2f_lw_RID               => hps_h2f_lw_axi_master_rid,       --                  .rid
			h2f_lw_RDATA             => hps_h2f_lw_axi_master_rdata,     --                  .rdata
			h2f_lw_RRESP             => hps_h2f_lw_axi_master_rresp,     --                  .rresp
			h2f_lw_RLAST             => hps_h2f_lw_axi_master_rlast,     --                  .rlast
			h2f_lw_RVALID            => hps_h2f_lw_axi_master_rvalid,    --                  .rvalid
			h2f_lw_RREADY            => hps_h2f_lw_axi_master_rready,    --                  .rready
			f2h_irq_p0               => hps_f2h_irq0_irq,                --          f2h_irq0.irq
			f2h_irq_p1               => hps_f2h_irq1_irq                 --          f2h_irq1.irq
		);

	led : component soc_system_led
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => led_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => led_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => led_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => led_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => led_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => led_external_connection_export                         -- external_connection.export
		);

	pb : component soc_system_pb
		port map (
			clk      => clk_clk,                                       --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => pb_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => pb_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => pb_external_connection_export                  -- external_connection.export
		);

	lfsr_0 : component number_generator
		port map (
			reset_in => rst_controller_reset_out_reset_ports_inv,                        --          reset.reset_n
			clk_in   => clk_clk,                                                         --          clock.clk
			CS       => lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect, -- avalon_slave_0.chipselect
			OE       => lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_read,       --               .read
			readdata => lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata    --               .readdata
		);

	led_s1_translator : component soc_system_led_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                    reset.reset
			uav_address              => led_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => led_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => led_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => led_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => led_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => led_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => led_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => led_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => led_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => led_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => led_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	pb_s1_translator : component soc_system_pb_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                   --                    reset.reset
			uav_address              => pb_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pb_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pb_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pb_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pb_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pb_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pb_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pb_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pb_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pb_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pb_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pb_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => pb_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                             --              (terminated)
			av_read                  => open,                                                             --              (terminated)
			av_writedata             => open,                                                             --              (terminated)
			av_begintransfer         => open,                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                             --              (terminated)
			av_burstcount            => open,                                                             --              (terminated)
			av_byteenable            => open,                                                             --              (terminated)
			av_readdatavalid         => '0',                                                              --              (terminated)
			av_waitrequest           => '0',                                                              --              (terminated)
			av_writebyteenable       => open,                                                             --              (terminated)
			av_lock                  => open,                                                             --              (terminated)
			av_chipselect            => open,                                                             --              (terminated)
			av_clken                 => open,                                                             --              (terminated)
			uav_clken                => '0',                                                              --              (terminated)
			av_debugaccess           => open,                                                             --              (terminated)
			av_outputenable          => open,                                                             --              (terminated)
			uav_response             => open,                                                             --              (terminated)
			av_response              => "00",                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                             --              (terminated)
			av_writeresponserequest  => open,                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                               --              (terminated)
		);

	lfsr_0_avalon_slave_0_translator : component soc_system_lfsr_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_read                  => lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --      avalon_anti_slave_0.read
			av_readdata              => lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_chipselect            => lfsr_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_address               => open,                                                                             --              (terminated)
			av_write                 => open,                                                                             --              (terminated)
			av_writedata             => open,                                                                             --              (terminated)
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_byteenable            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_debugaccess           => open,                                                                             --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	hps_h2f_lw_axi_master_agent : component altera_merlin_axi_master_ni
		generic map (
			ID_WIDTH                  => 12,
			ADDR_WIDTH                => 21,
			RDATA_WIDTH               => 32,
			WDATA_WIDTH               => 32,
			ADDR_USER_WIDTH           => 1,
			DATA_USER_WIDTH           => 1,
			AXI_BURST_LENGTH_WIDTH    => 4,
			AXI_LOCK_WIDTH            => 2,
			AXI_VERSION               => "AXI3",
			WRITE_ISSUING_CAPABILITY  => 8,
			READ_ISSUING_CAPABILITY   => 8,
			PKT_BEGIN_BURST           => 84,
			PKT_CACHE_H               => 108,
			PKT_CACHE_L               => 105,
			PKT_ADDR_SIDEBAND_H       => 82,
			PKT_ADDR_SIDEBAND_L       => 82,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_EXCLUSIVE       => 62,
			PKT_TRANS_LOCK            => 61,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 101,
			PKT_THREAD_ID_L           => 90,
			PKT_QOS_L                 => 85,
			PKT_QOS_H                 => 85,
			PKT_DATA_SIDEBAND_H       => 83,
			PKT_DATA_SIDEBAND_L       => 83,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 3,
			ID                        => 0
		)
		port map (
			aclk                   => clk_clk,                                            --              clk.clk
			aresetn                => rst_controller_reset_out_reset_ports_inv,           --        clk_reset.reset_n
			write_cp_valid         => hps_h2f_lw_axi_master_agent_write_cp_valid,         --         write_cp.valid
			write_cp_data          => hps_h2f_lw_axi_master_agent_write_cp_data,          --                 .data
			write_cp_startofpacket => hps_h2f_lw_axi_master_agent_write_cp_startofpacket, --                 .startofpacket
			write_cp_endofpacket   => hps_h2f_lw_axi_master_agent_write_cp_endofpacket,   --                 .endofpacket
			write_cp_ready         => hps_h2f_lw_axi_master_agent_write_cp_ready,         --                 .ready
			write_rp_valid         => limiter_rsp_src_valid,                              --         write_rp.valid
			write_rp_data          => limiter_rsp_src_data,                               --                 .data
			write_rp_channel       => limiter_rsp_src_channel,                            --                 .channel
			write_rp_startofpacket => limiter_rsp_src_startofpacket,                      --                 .startofpacket
			write_rp_endofpacket   => limiter_rsp_src_endofpacket,                        --                 .endofpacket
			write_rp_ready         => limiter_rsp_src_ready,                              --                 .ready
			read_cp_valid          => hps_h2f_lw_axi_master_agent_read_cp_valid,          --          read_cp.valid
			read_cp_data           => hps_h2f_lw_axi_master_agent_read_cp_data,           --                 .data
			read_cp_startofpacket  => hps_h2f_lw_axi_master_agent_read_cp_startofpacket,  --                 .startofpacket
			read_cp_endofpacket    => hps_h2f_lw_axi_master_agent_read_cp_endofpacket,    --                 .endofpacket
			read_cp_ready          => hps_h2f_lw_axi_master_agent_read_cp_ready,          --                 .ready
			read_rp_valid          => limiter_001_rsp_src_valid,                          --          read_rp.valid
			read_rp_data           => limiter_001_rsp_src_data,                           --                 .data
			read_rp_channel        => limiter_001_rsp_src_channel,                        --                 .channel
			read_rp_startofpacket  => limiter_001_rsp_src_startofpacket,                  --                 .startofpacket
			read_rp_endofpacket    => limiter_001_rsp_src_endofpacket,                    --                 .endofpacket
			read_rp_ready          => limiter_001_rsp_src_ready,                          --                 .ready
			awid                   => hps_h2f_lw_axi_master_awid,                         -- altera_axi_slave.awid
			awaddr                 => hps_h2f_lw_axi_master_awaddr,                       --                 .awaddr
			awlen                  => hps_h2f_lw_axi_master_awlen,                        --                 .awlen
			awsize                 => hps_h2f_lw_axi_master_awsize,                       --                 .awsize
			awburst                => hps_h2f_lw_axi_master_awburst,                      --                 .awburst
			awlock                 => hps_h2f_lw_axi_master_awlock,                       --                 .awlock
			awcache                => hps_h2f_lw_axi_master_awcache,                      --                 .awcache
			awprot                 => hps_h2f_lw_axi_master_awprot,                       --                 .awprot
			awvalid                => hps_h2f_lw_axi_master_awvalid,                      --                 .awvalid
			awready                => hps_h2f_lw_axi_master_awready,                      --                 .awready
			wid                    => hps_h2f_lw_axi_master_wid,                          --                 .wid
			wdata                  => hps_h2f_lw_axi_master_wdata,                        --                 .wdata
			wstrb                  => hps_h2f_lw_axi_master_wstrb,                        --                 .wstrb
			wlast                  => hps_h2f_lw_axi_master_wlast,                        --                 .wlast
			wvalid                 => hps_h2f_lw_axi_master_wvalid,                       --                 .wvalid
			wready                 => hps_h2f_lw_axi_master_wready,                       --                 .wready
			bid                    => hps_h2f_lw_axi_master_bid,                          --                 .bid
			bresp                  => hps_h2f_lw_axi_master_bresp,                        --                 .bresp
			bvalid                 => hps_h2f_lw_axi_master_bvalid,                       --                 .bvalid
			bready                 => hps_h2f_lw_axi_master_bready,                       --                 .bready
			arid                   => hps_h2f_lw_axi_master_arid,                         --                 .arid
			araddr                 => hps_h2f_lw_axi_master_araddr,                       --                 .araddr
			arlen                  => hps_h2f_lw_axi_master_arlen,                        --                 .arlen
			arsize                 => hps_h2f_lw_axi_master_arsize,                       --                 .arsize
			arburst                => hps_h2f_lw_axi_master_arburst,                      --                 .arburst
			arlock                 => hps_h2f_lw_axi_master_arlock,                       --                 .arlock
			arcache                => hps_h2f_lw_axi_master_arcache,                      --                 .arcache
			arprot                 => hps_h2f_lw_axi_master_arprot,                       --                 .arprot
			arvalid                => hps_h2f_lw_axi_master_arvalid,                      --                 .arvalid
			arready                => hps_h2f_lw_axi_master_arready,                      --                 .arready
			rid                    => hps_h2f_lw_axi_master_rid,                          --                 .rid
			rdata                  => hps_h2f_lw_axi_master_rdata,                        --                 .rdata
			rresp                  => hps_h2f_lw_axi_master_rresp,                        --                 .rresp
			rlast                  => hps_h2f_lw_axi_master_rlast,                        --                 .rlast
			rvalid                 => hps_h2f_lw_axi_master_rvalid,                       --                 .rvalid
			rready                 => hps_h2f_lw_axi_master_rready,                       --                 .rready
			awuser                 => "0",                                                --      (terminated)
			aruser                 => "0",                                                --      (terminated)
			awqos                  => "0000",                                             --      (terminated)
			arqos                  => "0000",                                             --      (terminated)
			awregion               => "0000",                                             --      (terminated)
			arregion               => "0000",                                             --      (terminated)
			wuser                  => "0",                                                --      (terminated)
			ruser                  => open,                                               --      (terminated)
			buser                  => open                                                --      (terminated)
		);

	led_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 3,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => led_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => led_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => led_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => led_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => led_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => led_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => led_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => led_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => led_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                 --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                 --                .valid
			cp_data                 => burst_adapter_source0_data,                                                  --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                           --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                               --                .channel
			rf_sink_ready           => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 112,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			in_data           => led_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			in_data           => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                  -- (terminated)
			csr_read          => '0',                                                                   -- (terminated)
			csr_write         => '0',                                                                   -- (terminated)
			csr_readdata      => open,                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                    -- (terminated)
			almost_full_data  => open,                                                                  -- (terminated)
			almost_empty_data => open,                                                                  -- (terminated)
			in_startofpacket  => '0',                                                                   -- (terminated)
			in_endofpacket    => '0',                                                                   -- (terminated)
			out_startofpacket => open,                                                                  -- (terminated)
			out_endofpacket   => open,                                                                  -- (terminated)
			in_empty          => '0',                                                                   -- (terminated)
			out_empty         => open,                                                                  -- (terminated)
			in_error          => '0',                                                                   -- (terminated)
			out_error         => open,                                                                  -- (terminated)
			in_channel        => '0',                                                                   -- (terminated)
			out_channel       => open                                                                   -- (terminated)
		);

	pb_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 3,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                             --       clk_reset.reset
			m0_address              => pb_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pb_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pb_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pb_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pb_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pb_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pb_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pb_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pb_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pb_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pb_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pb_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pb_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pb_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pb_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pb_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                            --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                            --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                             --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                    --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                      --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                          --                .channel
			rf_sink_ready           => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                         --     (terminated)
		);

	pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 112,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                             -- clk_reset.reset
			in_data           => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pb_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pb_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                       -- (terminated)
			csr_read          => '0',                                                                        -- (terminated)
			csr_write         => '0',                                                                        -- (terminated)
			csr_readdata      => open,                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                         -- (terminated)
			almost_full_data  => open,                                                                       -- (terminated)
			almost_empty_data => open,                                                                       -- (terminated)
			in_empty          => '0',                                                                        -- (terminated)
			out_empty         => open,                                                                       -- (terminated)
			in_error          => '0',                                                                        -- (terminated)
			out_error         => open,                                                                       -- (terminated)
			in_channel        => '0',                                                                        -- (terminated)
			out_channel       => open                                                                        -- (terminated)
		);

	pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			in_data           => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => pb_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                 -- (terminated)
			csr_read          => '0',                                                                  -- (terminated)
			csr_write         => '0',                                                                  -- (terminated)
			csr_readdata      => open,                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                   -- (terminated)
			almost_full_data  => open,                                                                 -- (terminated)
			almost_empty_data => open,                                                                 -- (terminated)
			in_startofpacket  => '0',                                                                  -- (terminated)
			in_endofpacket    => '0',                                                                  -- (terminated)
			out_startofpacket => open,                                                                 -- (terminated)
			out_endofpacket   => open,                                                                 -- (terminated)
			in_empty          => '0',                                                                  -- (terminated)
			out_empty         => open,                                                                 -- (terminated)
			in_error          => '0',                                                                  -- (terminated)
			out_error         => open,                                                                 -- (terminated)
			in_channel        => '0',                                                                  -- (terminated)
			out_channel       => open                                                                  -- (terminated)
		);

	lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 3,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_002_source0_ready,                                                            --              cp.ready
			cp_valid                => burst_adapter_002_source0_valid,                                                            --                .valid
			cp_data                 => burst_adapter_002_source0_data,                                                             --                .data
			cp_startofpacket        => burst_adapter_002_source0_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => burst_adapter_002_source0_endofpacket,                                                      --                .endofpacket
			cp_channel              => burst_adapter_002_source0_channel,                                                          --                .channel
			rf_sink_ready           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 112,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo : component soc_system_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                 -- (terminated)
			csr_read          => '0',                                                                                  -- (terminated)
			csr_write         => '0',                                                                                  -- (terminated)
			csr_readdata      => open,                                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                   -- (terminated)
			almost_full_data  => open,                                                                                 -- (terminated)
			almost_empty_data => open,                                                                                 -- (terminated)
			in_startofpacket  => '0',                                                                                  -- (terminated)
			in_endofpacket    => '0',                                                                                  -- (terminated)
			out_startofpacket => open,                                                                                 -- (terminated)
			out_endofpacket   => open,                                                                                 -- (terminated)
			in_empty          => '0',                                                                                  -- (terminated)
			out_empty         => open,                                                                                 -- (terminated)
			in_error          => '0',                                                                                  -- (terminated)
			out_error         => open,                                                                                 -- (terminated)
			in_channel        => '0',                                                                                  -- (terminated)
			out_channel       => open                                                                                  -- (terminated)
		);

	addr_router : component soc_system_addr_router
		port map (
			sink_ready         => hps_h2f_lw_axi_master_agent_write_cp_ready,         --      sink.ready
			sink_valid         => hps_h2f_lw_axi_master_agent_write_cp_valid,         --          .valid
			sink_data          => hps_h2f_lw_axi_master_agent_write_cp_data,          --          .data
			sink_startofpacket => hps_h2f_lw_axi_master_agent_write_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => hps_h2f_lw_axi_master_agent_write_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                              --       src.ready
			src_valid          => addr_router_src_valid,                              --          .valid
			src_data           => addr_router_src_data,                               --          .data
			src_channel        => addr_router_src_channel,                            --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                      --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                         --          .endofpacket
		);

	addr_router_001 : component soc_system_addr_router
		port map (
			sink_ready         => hps_h2f_lw_axi_master_agent_read_cp_ready,         --      sink.ready
			sink_valid         => hps_h2f_lw_axi_master_agent_read_cp_valid,         --          .valid
			sink_data          => hps_h2f_lw_axi_master_agent_read_cp_data,          --          .data
			sink_startofpacket => hps_h2f_lw_axi_master_agent_read_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => hps_h2f_lw_axi_master_agent_read_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                    -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                         --       src.ready
			src_valid          => addr_router_001_src_valid,                         --          .valid
			src_data           => addr_router_001_src_data,                          --          .data
			src_channel        => addr_router_001_src_channel,                       --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                 --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                    --          .endofpacket
		);

	id_router : component soc_system_id_router
		port map (
			sink_ready         => led_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => led_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => led_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_src_ready,                                               --       src.ready
			src_valid          => id_router_src_valid,                                               --          .valid
			src_data           => id_router_src_data,                                                --          .data
			src_channel        => id_router_src_channel,                                             --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                          --          .endofpacket
		);

	id_router_001 : component soc_system_id_router
		port map (
			sink_ready         => pb_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pb_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pb_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pb_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pb_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                   -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                          --       src.ready
			src_valid          => id_router_001_src_valid,                                          --          .valid
			src_data           => id_router_001_src_data,                                           --          .data
			src_channel        => id_router_001_src_channel,                                        --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                  --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                     --          .endofpacket
		);

	id_router_002 : component soc_system_id_router
		port map (
			sink_ready         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lfsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                          --       src.ready
			src_valid          => id_router_002_src_valid,                                                          --          .valid
			src_data           => id_router_002_src_data,                                                           --          .data
			src_channel        => id_router_002_src_channel,                                                        --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                     --          .endofpacket
		);

	limiter : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			MAX_OUTSTANDING_RESPONSES => 3,
			PIPELINED                 => 0,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 3,
			VALID_WIDTH               => 3,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_clk,                        --       clk.clk
			reset                  => rst_controller_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,          --          .valid
			cmd_sink_data          => addr_router_src_data,           --          .data
			cmd_sink_channel       => addr_router_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data          -- cmd_valid.data
		);

	limiter_001 : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			MAX_OUTSTANDING_RESPONSES => 3,
			PIPELINED                 => 0,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 3,
			VALID_WIDTH               => 3,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_clk,                            --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_001_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_001_src_valid,          --          .valid
			cmd_sink_data          => addr_router_001_src_data,           --          .data
			cmd_sink_channel       => addr_router_001_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_001_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_001_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_001_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_001_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_001_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_001_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_001_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_001_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_001_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_001_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_001_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_001_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_001_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_001_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_001_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_001_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_001_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_001_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_001_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_001_cmd_valid_data          -- cmd_valid.data
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_BEGIN_BURST           => 84,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 70,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 1,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 3,
			OUT_BYTE_CNT_H            => 65,
			OUT_BURSTWRAP_H           => 76,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 0,
			BURSTWRAP_CONST_VALUE     => 0
		)
		port map (
			clk                   => clk_clk,                             --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_src_ready,              --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_BEGIN_BURST           => 84,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 70,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 1,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 3,
			OUT_BYTE_CNT_H            => 65,
			OUT_BURSTWRAP_H           => 76,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 0,
			BURSTWRAP_CONST_VALUE     => 0
		)
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_001_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_001_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_001_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_001_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_001_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_001_src_ready,              --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	burst_adapter_002 : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_BEGIN_BURST           => 84,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 63,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 70,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 1,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 3,
			OUT_BYTE_CNT_H            => 65,
			OUT_BURSTWRAP_H           => 76,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 0,
			BURSTWRAP_CONST_VALUE     => 0
		)
		port map (
			clk                   => clk_clk,                                 --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_002_src_valid,              --     sink0.valid
			sink0_data            => cmd_xbar_mux_002_src_data,               --          .data
			sink0_channel         => cmd_xbar_mux_002_src_channel,            --          .channel
			sink0_startofpacket   => cmd_xbar_mux_002_src_startofpacket,      --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_002_src_endofpacket,        --          .endofpacket
			sink0_ready           => cmd_xbar_mux_002_src_ready,              --          .ready
			source0_valid         => burst_adapter_002_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_002_source0_data,          --          .data
			source0_channel       => burst_adapter_002_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_002_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_002_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_002_source0_ready          --          .ready
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => hps_h2f_reset_reset_ports_inv,  -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	cmd_xbar_demux : component soc_system_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --        clk.clk
			reset              => rst_controller_reset_out_reset,    --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_cmd_src_channel,           --           .channel
			sink_data          => limiter_cmd_src_data,              --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_001 : component soc_system_cmd_xbar_demux
		port map (
			clk                => clk_clk,                               --        clk.clk
			reset              => rst_controller_reset_out_reset,        --  clk_reset.reset
			sink_ready         => limiter_001_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_001_cmd_src_channel,           --           .channel
			sink_data          => limiter_001_cmd_src_data,              --           .data
			sink_startofpacket => limiter_001_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_001_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_001_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --           .endofpacket
		);

	cmd_xbar_mux : component soc_system_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component soc_system_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component soc_system_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component soc_system_rsp_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component soc_system_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component soc_system_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component soc_system_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component soc_system_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk        => open,             --       clk.clk
			reset      => open,             -- clk_reset.reset
			sender_irq => hps_f2h_irq0_irq  --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper
		port map (
			clk        => open,             --       clk.clk
			reset      => open,             -- clk_reset.reset
			sender_irq => hps_f2h_irq1_irq  --    sender.irq
		);

	led_s1_translator_avalon_anti_slave_0_write_ports_inv <= not led_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_h2f_reset_reset_ports_inv <= not hps_h2f_reset_reset;

end architecture rtl; -- of soc_system
