-- megafunction wizard: %FIR Compiler II v13.0%
-- GENERATION: XML
-- fir.vhd

-- Generated using ACDS version 13.0sp1 232 at 2016.05.11.17:50:50

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fir is
	port (
		clk              : in  std_logic                     := '0';             --                     clk.clk
		reset_n          : in  std_logic                     := '0';             --                     rst.reset_n
		ast_sink_data    : in  std_logic_vector(16 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                     := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(36 downto 0);                    -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                        --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0)                      --                        .error
	);
end entity fir;

architecture rtl of fir is
	component fir_0002 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(16 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(36 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                      -- error
		);
	end component fir_0002;

begin

	fir_inst : component fir_0002
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of fir
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.0" >
-- Retrieval info: 	<generic name="deviceFamily" value="Cyclone V" />
-- Retrieval info: 	<generic name="filterType" value="Single Rate" />
-- Retrieval info: 	<generic name="interpFactor" value="1" />
-- Retrieval info: 	<generic name="decimFactor" value="1" />
-- Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
-- Retrieval info: 	<generic name="clockRate" value="65" />
-- Retrieval info: 	<generic name="clockSlack" value="0" />
-- Retrieval info: 	<generic name="speedGrade" value="Medium" />
-- Retrieval info: 	<generic name="coeffReload" value="false" />
-- Retrieval info: 	<generic name="baseAddress" value="0" />
-- Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
-- Retrieval info: 	<generic name="backPressure" value="false" />
-- Retrieval info: 	<generic name="symmetryMode" value="Non Symmetry" />
-- Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
-- Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
-- Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
-- Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
-- Retrieval info: 	<generic name="inputRate" value="65" />
-- Retrieval info: 	<generic name="inputChannelNum" value="1" />
-- Retrieval info: 	<generic name="inputType" value="Signed Binary" />
-- Retrieval info: 	<generic name="inputBitWidth" value="14" />
-- Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffSetRealValue" value="0.007587141,-0.00712971,-0.005379073,-0.004540912,-0.004147896,-0.003910773,-0.003665469,-0.00330336,-0.002767768,-0.002036356,-0.001114017,-2.452896E-5,0.001186563,0.002457356,0.003712499,0.00487123,0.005848455,0.00656088,0.006930976,0.006896451,0.006413709,0.005463123,0.00404986,0.002209181,6.840301E-6,-0.002460025,-0.005068684,-0.007674145,-0.01011588,-0.01222235,-0.01382094,-0.01474603,-0.01484945,-0.01400697,-0.01212771,-0.009161554,-0.005106092,-6.874279E-6,0.006044521,0.01291255,0.02041769,0.02833927,0.03642753,0.04441774,0.05204455,0.0590423,0.06515768,0.07015625,0.07387265,0.07616962,0.07692465,0.07616962,0.07387265,0.07015625,0.06515768,0.0590423,0.05204455,0.04441774,0.03642753,0.02833927,0.02041769,0.01291255,0.006044521,-6.874279E-6,-0.005106092,-0.009161554,-0.01212771,-0.01400697,-0.01484945,-0.01474603,-0.01382094,-0.01222235,-0.01011588,-0.007674145,-0.005068684,-0.002460025,6.840301E-6,0.002209181,0.00404986,0.005463123,0.006413709,0.006896451,0.006930976,0.00656088,0.005848455,0.00487123,0.003712499,0.002457356,0.001186563,-2.452896E-5,-0.001114017,-0.002036356,-0.002767768,-0.00330336,-0.003665469,-0.003910773,-0.004147896,-0.004540912,-0.005379073,-0.00712971,0.007587141,-0.00657841,0.008071934,0.005793007,0.004662922,0.0037703,0.002677979,0.001253782,-4.294037E-4,-0.002140719,-0.003584093,-0.004458208,-0.004528231,-0.003691834,-0.002014937,2.618153E-4,0.002752052,0.004980554,0.006468821,0.006835354,0.005878667,0.003637662,4.096352E-4,-0.003276936,-0.006741182,-0.009268469,-0.01024592,-0.009293643,-0.006364493,-0.001791119,0.003730613,0.009231984,0.01362203,0.01588133,0.01526181,0.01145918,0.004729703,-0.004081433,-0.01360557,-0.02211112,-0.02774294,-0.02880796,-0.02406421,-0.0129438,0.004304452,0.02656958,0.05196313,0.07802749,0.1020776,0.1215001,0.1340984,0.138483,0.1340984,0.1215001,0.1020776,0.07802749,0.05196313,0.02656958,0.004304452,-0.0129438,-0.02406421,-0.02880796,-0.02774294,-0.02211112,-0.01360557,-0.004081433,0.004729703,0.01145918,0.01526181,0.01588133,0.01362203,0.009231984,0.003730613,-0.001791119,-0.006364493,-0.009293643,-0.01024592,-0.009268469,-0.006741182,-0.003276936,4.096352E-4,0.003637662,0.005878667,0.006835354,0.006468821,0.004980554,0.002752052,2.618153E-4,-0.002014937,-0.003691834,-0.004528231,-0.004458208,-0.003584093,-0.002140719,-4.294037E-4,0.001253782,0.002677979,0.0037703,0.004662922,0.005793007,0.008071934,-0.00657841,-0.007587141,0.00712971,0.005379073,0.004540912,0.004147896,0.003910773,0.003665469,0.00330336,0.002767768,0.002036356,0.001114017,2.452896E-5,-0.001186563,-0.002457356,-0.003712499,-0.00487123,-0.005848455,-0.00656088,-0.006930976,-0.006896451,-0.006413709,-0.005463123,-0.00404986,-0.002209181,-6.840301E-6,0.002460025,0.005068684,0.007674145,0.01011588,0.01222235,0.01382094,0.01474603,0.01484945,0.01400697,0.01212771,0.009161554,0.005106092,6.874279E-6,-0.006044521,-0.01291255,-0.02041769,-0.02833927,-0.03642753,-0.04441774,-0.05204455,-0.0590423,-0.06515768,-0.07015625,-0.07387265,-0.07616962,0.9230754,-0.07616962,-0.07387265,-0.07015625,-0.06515768,-0.0590423,-0.05204455,-0.04441774,-0.03642753,-0.02833927,-0.02041769,-0.01291255,-0.006044521,6.874279E-6,0.005106092,0.009161554,0.01212771,0.01400697,0.01484945,0.01474603,0.01382094,0.01222235,0.01011588,0.007674145,0.005068684,0.002460025,-6.840301E-6,-0.002209181,-0.00404986,-0.005463123,-0.006413709,-0.006896451,-0.006930976,-0.00656088,-0.005848455,-0.00487123,-0.003712499,-0.002457356,-0.001186563,2.452896E-5,0.001114017,0.002036356,0.002767768,0.00330336,0.003665469,0.003910773,0.004147896,0.004540912,0.005379073,0.00712971,-0.007587141,0.00657841,-0.008071934,-0.005793007,-0.004662922,-0.0037703,-0.002677979,-0.001253782,4.294037E-4,0.002140719,0.003584093,0.004458208,0.004528231,0.003691834,0.002014937,-2.618153E-4,-0.002752052,-0.004980554,-0.006468821,-0.006835354,-0.005878667,-0.003637662,-4.096352E-4,0.003276936,0.006741182,0.009268469,0.01024592,0.009293643,0.006364493,0.001791119,-0.003730613,-0.009231984,-0.01362203,-0.01588133,-0.01526181,-0.01145918,-0.004729703,0.004081433,0.01360557,0.02211112,0.02774294,0.02880796,0.02406421,0.0129438,-0.004304452,-0.02656958,-0.05196313,-0.07802749,-0.1020776,-0.1215001,-0.1340984,0.861517,-0.1340984,-0.1215001,-0.1020776,-0.07802749,-0.05196313,-0.02656958,-0.004304452,0.0129438,0.02406421,0.02880796,0.02774294,0.02211112,0.01360557,0.004081433,-0.004729703,-0.01145918,-0.01526181,-0.01588133,-0.01362203,-0.009231984,-0.003730613,0.001791119,0.006364493,0.009293643,0.01024592,0.009268469,0.006741182,0.003276936,-4.096352E-4,-0.003637662,-0.005878667,-0.006835354,-0.006468821,-0.004980554,-0.002752052,-2.618153E-4,0.002014937,0.003691834,0.004528231,0.004458208,0.003584093,0.002140719,4.294037E-4,-0.001253782,-0.002677979,-0.0037703,-0.004662922,-0.005793007,-0.008071934,0.00657841,-0.01535534,0.003844121,0.003356547,0.002812384,0.002129428,0.001257891,2.237009E-4,-8.67154E-4,-0.001825938,-0.002421135,-0.002408962,-0.001606216,6.238768E-5,0.002506686,0.0054929,0.008633849,0.01144432,0.01344879,0.01423409,0.0135682,0.01144893,0.0081365,0.00412478,7.108923E-5,-0.003313962,-0.005407756,-0.005803749,-0.004424986,-0.00156611,0.00209793,0.00561796,0.007910996,0.007944382,0.004956525,-0.001372941,-0.01079768,-0.02246449,-0.03497623,-0.04655265,-0.0552799,-0.05938353,-0.05753765,-0.04907087,-0.03421436,-0.01398309,0.009719415,0.03444171,0.05749471,0.07623178,0.08845544,0.09269743,0.08845544,0.07623178,0.05749471,0.03444171,0.009719415,-0.01398309,-0.03421436,-0.04907087,-0.05753765,-0.05938353,-0.0552799,-0.04655265,-0.03497623,-0.02246449,-0.01079768,-0.001372941,0.004956525,0.007944382,0.007910996,0.00561796,0.00209793,-0.00156611,-0.004424986,-0.005803749,-0.005407756,-0.003313962,7.108923E-5,0.00412478,0.0081365,0.01144893,0.0135682,0.01423409,0.01344879,0.01144432,0.008633849,0.0054929,0.002506686,6.238768E-5,-0.001606216,-0.002408962,-0.002421135,-0.001825938,-8.67154E-4,2.237009E-4,0.001257891,0.002129428,0.002812384,0.003356547,0.003844121,-0.01535534,0.004771988,-0.004521916,0.007701157,0.005817928,-0.001461344,-0.006927878,-0.00858482,-0.007255783,-0.00436718,-0.001434061,3.902571E-5,-7.136291E-4,-0.002979765,-0.004685495,-0.003636287,8.846245E-4,0.007275901,0.01232731,0.01306836,0.008726895,0.001439445,-0.004875604,-0.006964929,-0.004379524,9.374849E-6,0.001730203,-0.002235362,-0.01104012,-0.01990814,-0.02267321,-0.01573227,-7.576433E-4,0.01560104,0.02530153,0.02389398,0.01363022,0.002656234,2.537939E-5,0.009497112,0.02578941,0.03622342,0.02758404,-0.005255461,-0.05392099,-0.09816467,-0.1146139,-0.08871266,-0.02362953,0.05895042,0.1273164,0.1537509,0.1273164,0.05895042,-0.02362953,-0.08871266,-0.1146139,-0.09816467,-0.05392099,-0.005255461,0.02758404,0.03622342,0.02578941,0.009497112,2.537939E-5,0.002656234,0.01363022,0.02389398,0.02530153,0.01560104,-7.576433E-4,-0.01573227,-0.02267321,-0.01990814,-0.01104012,-0.002235362,0.001730203,9.374849E-6,-0.004379524,-0.006964929,-0.004875604,0.001439445,0.008726895,0.01306836,0.01232731,0.007275901,8.846245E-4,-0.003636287,-0.004685495,-0.002979765,-7.136291E-4,3.902571E-5,-0.001434061,-0.00436718,-0.007255783,-0.00858482,-0.006927878,-0.001461344,0.005817928,0.007701157,-0.004521916,0.004771988,0.01535534,-0.003844121,-0.003356547,-0.002812384,-0.002129428,-0.001257891,-2.237009E-4,8.67154E-4,0.001825938,0.002421135,0.002408962,0.001606216,-6.238768E-5,-0.002506686,-0.0054929,-0.008633849,-0.01144432,-0.01344879,-0.01423409,-0.0135682,-0.01144893,-0.0081365,-0.00412478,-7.108923E-5,0.003313962,0.005407756,0.005803749,0.004424986,0.00156611,-0.00209793,-0.00561796,-0.007910996,-0.007944382,-0.004956525,0.001372941,0.01079768,0.02246449,0.03497623,0.04655265,0.0552799,0.05938353,0.05753765,0.04907087,0.03421436,0.01398309,-0.009719415,-0.03444171,-0.05749471,-0.07623178,-0.08845544,0.9073026,-0.08845544,-0.07623178,-0.05749471,-0.03444171,-0.009719415,0.01398309,0.03421436,0.04907087,0.05753765,0.05938353,0.0552799,0.04655265,0.03497623,0.02246449,0.01079768,0.001372941,-0.004956525,-0.007944382,-0.007910996,-0.00561796,-0.00209793,0.00156611,0.004424986,0.005803749,0.005407756,0.003313962,-7.108923E-5,-0.00412478,-0.0081365,-0.01144893,-0.0135682,-0.01423409,-0.01344879,-0.01144432,-0.008633849,-0.0054929,-0.002506686,-6.238768E-5,0.001606216,0.002408962,0.002421135,0.001825938,8.67154E-4,-2.237009E-4,-0.001257891,-0.002129428,-0.002812384,-0.003356547,-0.003844121,0.01535534,-0.004771988,0.004521916,-0.007701157,-0.005817928,0.001461344,0.006927878,0.00858482,0.007255783,0.00436718,0.001434061,-3.902571E-5,7.136291E-4,0.002979765,0.004685495,0.003636287,-8.846245E-4,-0.007275901,-0.01232731,-0.01306836,-0.008726895,-0.001439445,0.004875604,0.006964929,0.004379524,-9.374849E-6,-0.001730203,0.002235362,0.01104012,0.01990814,0.02267321,0.01573227,7.576433E-4,-0.01560104,-0.02530153,-0.02389398,-0.01363022,-0.002656234,-2.537939E-5,-0.009497112,-0.02578941,-0.03622342,-0.02758404,0.005255461,0.05392099,0.09816467,0.1146139,0.08871266,0.02362953,-0.05895042,-0.1273164,0.8462491,-0.1273164,-0.05895042,0.02362953,0.08871266,0.1146139,0.09816467,0.05392099,0.005255461,-0.02758404,-0.03622342,-0.02578941,-0.009497112,-2.537939E-5,-0.002656234,-0.01363022,-0.02389398,-0.02530153,-0.01560104,7.576433E-4,0.01573227,0.02267321,0.01990814,0.01104012,0.002235362,-0.001730203,-9.374849E-6,0.004379524,0.006964929,0.004875604,-0.001439445,-0.008726895,-0.01306836,-0.01232731,-0.007275901,-8.846245E-4,0.003636287,0.004685495,0.002979765,7.136291E-4,-3.902571E-5,0.001434061,0.00436718,0.007255783,0.00858482,0.006927878,0.001461344,-0.005817928,-0.007701157,0.004521916,-0.004771988" />
-- Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
-- Retrieval info: 	<generic name="coeffScaling" value="Auto" />
-- Retrieval info: 	<generic name="coeffBitWidth" value="16" />
-- Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="outType" value="Signed Binary" />
-- Retrieval info: 	<generic name="outMSBRound" value="Truncation" />
-- Retrieval info: 	<generic name="outMsbBitRem" value="0" />
-- Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
-- Retrieval info: 	<generic name="outLsbBitRem" value="0" />
-- Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
-- Retrieval info: 	<generic name="bankCount" value="8" />
-- Retrieval info: 	<generic name="bankDisplay" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : NONE
